

module top (
    
);

endmodule
