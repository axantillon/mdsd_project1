/*
    Diego Bonilla, Enrique Macaya, Sebastian Lopez, Andres Antillon
    Project 1
    ECE 2372
    Dr. Juan Carlos Rojas
    Register module
*/


module alu(input OP[0:3], input A[0:7], input B[0:7], output Z[0:7]);

endmodule