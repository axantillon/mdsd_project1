/*
    Diego Bonilla, Enrique Macaya, Sebastian Lopez, Andres Antillon
    Project 1
    ECE 2372
    Dr. Juan Carlos Rojas
    Testbench
*/

module alu_testbench();

endmodule

module register_testbench();

endmodule

module datapath_testbench();

endmodule