

module instructionMemory (
    input wire [7:0] address,
    input wire [1:0] programSelect,
    output wire [15:0] instruction
);

    reg [15:0] sumIntegersProgram [0:127] = '{
        8'd0: 16'b0010000000000001,
        8'd1: 16'b0010000000000010,
        8'd2: 16'b0010000000000011,
        8'd3: 16'b0010000000000100,
        8'd4: 16'b0010000000000101,
        8'd5: 16'b0010000000000110,
        8'd6: 16'b0010000000000111,
        8'd7: 16'b0010000000001000
    };

    reg [15:0] squareOfNProgram [0:127] = '{
        8'd0: 16'b0010000000000001,
        8'd1: 16'b0010000000000010,
        8'd2: 16'b0010000000000011,
        8'd3: 16'b0010000000000100,
        8'd4: 16'b0010000000000101,
        8'd5: 16'b0010000000000110,
        8'd6: 16'b0010000000000111,
        8'd7: 16'b0010000000001000
    };

    reg [15:0] 3Program [0:127] = '{
        8'd0: 16'b0010000000000001,
        8'd1: 16'b0010000000000010,
        8'd2: 16'b0010000000000011,
        8'd3: 16'b0010000000000100,
        8'd4: 16'b0010000000000101,
        8'd5: 16'b0010000000000110,
        8'd6: 16'b0010000000000111,
        8'd7: 16'b0010000000001000
    };

    reg [15:0] 4Program [0:127] = '{
        8'd0: 16'b0010000000000001,
        8'd1: 16'b0010000000000010,
        8'd2: 16'b0010000000000011,
        8'd3: 16'b0010000000000100,
        8'd4: 16'b0010000000000101,
        8'd5: 16'b0010000000000110,
        8'd6: 16'b0010000000000111,
        8'd7: 16'b0010000000001000
    };

    assign instruction =    programSelect == 2'b00 ? sumIntegersProgram[address] :
                            programSelect == 2'b01 ? squareOfNProgram[address] :
                            programSelect == 2'b10 ? 3Program[address] :
                            programSelect == 2'b11 ? 4Program[address] : 16'b0;

endmodule